LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all; 

ENTITY BF IS

PORT ( CLK, ENABLE: IN std_logic;
       AI,AR,BI,BR,WR,WI: IN SIGNED(19 downto 0); -- va cambiato il formato e conversioni
      SEL_INV,SEL3,SEL1,SELSUM,C,A_S,EN_REGR : IN std_logic;
		SEL2 : IN std_logic_vector(1 downto 0);
		EN_REGO : IN std_logic_vector(2 downto 0);
		A1R,A1I,B1R,B1I,AI_CTRL,AR_CTRL,BI_CTRL,BR_CTRL: OUT SIGNED(19 downto 0));
END BF;

ARCHITECTURE BEHAV OF BF IS 

COMPONENT RF IS
PORT ( CLK, ENABLE: IN std_logic;
       AI,AR,BI,BR,WR,WI: IN SIGNED(19 downto 0); -- va cambiato il formato e conversioni
      SEL3,SEL1 : IN std_logic;
		SEL2 : IN std_logic_vector(1 downto 0);
		OUT_MUX1,OUT_MUX2,OUT_MUX3,AI_CTRL,AR_CTRL,BI_CTRL,BR_CTRL: OUT SIGNED(19 downto 0));
END COMPONENT;


COMPONENT MOL IS
PORT ( C,CLK: IN std_logic;
       ADD1,ADD2: IN SIGNED(19 downto 0);
       RESULT: OUT SIGNED(38 downto 0));
END COMPONENT;

COMPONENT SUM IS
PORT ( A_S,CLK: IN std_logic;
       T1,T2: IN SIGNED(38 downto 0);
       RESULT: OUT SIGNED(39 downto 0));
END COMPONENT;

COMPONENT REG_39_M IS
PORT ( CLK: IN std_logic;
       D: IN SIGNED(38 downto 0);
       Q: OUT SIGNED(38 downto 0));
END COMPONENT;

COMPONENT REG_40_S IS
PORT ( CLK: IN std_logic;
       D: IN SIGNED(39 downto 0);
       Q: OUT SIGNED(39 downto 0));
END COMPONENT;

COMPONENT REG_ROUND IS
PORT ( CLK: IN std_logic;
		 ENABLE: IN std_logic;
       D: IN SIGNED(39 downto 0);
       Q: OUT SIGNED(39 downto 0));
END COMPONENT;

COMPONENT MUX39SUM IS 
PORT( A: IN SIGNED (19 downto 0); 			
		B: IN SIGNED(38 downto 0);				
		SEL : IN std_logic;
		OUTPUT: OUT SIGNED(38 downto 0));
END COMPONENT;

COMPONENT REG_A1R IS
PORT ( CLK: IN std_logic;
		 ENABLE: IN std_logic_vector(2 downto 0);
       D: IN SIGNED(19 downto 0);
       Q: OUT SIGNED(19 downto 0));
END COMPONENT;

COMPONENT REG_A1I IS
PORT ( CLK: IN std_logic;
		 ENABLE: IN std_logic_vector(2 downto 0);
       D: IN SIGNED(19 downto 0);
       Q: OUT SIGNED(19 downto 0));
END COMPONENT;

COMPONENT REG_B1R IS
PORT ( CLK: IN std_logic;
		 ENABLE: IN std_logic_vector(2 downto 0);
       D: IN SIGNED(19 downto 0);
       Q: OUT SIGNED(19 downto 0));
END COMPONENT;

COMPONENT REG_B1I IS
PORT ( CLK: IN std_logic;
		 ENABLE: IN std_logic_vector(2 downto 0);
       D: IN SIGNED(19 downto 0);
       Q: OUT SIGNED(19 downto 0));
END COMPONENT;

COMPONENT ROUNDING IS
PORT ( IN_39: IN SIGNED(39 downto 0);
       OUT_20: OUT SIGNED(19 downto 0));
END COMPONENT;

COMPONENT MUX_INV IS
PORT( A: IN SIGNED (38 downto 0);
		B: IN SIGNED(38 downto 0);
		SEL : IN std_logic;
		OUTPUT: OUT SIGNED(38 downto 0));
END COMPONENT;


SIGNAL BUSW,BUS1,BUS2,ROUNDED: SIGNED (19 downto 0);
SIGNAL MUXSUM_OUT,MOL_RES_IN,MOL_RES_OUT,OUTMUXINVT1,OUTMUXINVT2: SIGNED(38 downto 0);
SIGNAL SUM_RES_IN,SUM_RES_OUT,REG_ROUND_OUT: SIGNED(39 DOWNTO 0);
SIGNAL NOTHING: std_logic;
BEGIN 

ROUND: ROUNDING PORT MAP(IN_39=>REG_ROUND_OUT,OUT_20=>ROUNDED);
MUXSUM: MUX39SUM PORT MAP(A=>BUS1,B=>SUM_RES_OUT(38 DOWNTO 0),SEL=>SELSUM,OUTPUT=>MUXSUM_OUT);
REG_RF: RF PORT MAP (CLK=>CLK,ENABLE=>ENABLE,AI=>AI,AR=>AR,BI=>BI,BR=>BR,WR=>WR,WI=>WI,
							SEL1=>SEL1,SEL2=>SEL2,SEL3=>SEL3,AI_CTRL=>AI_CTRL,AR_CTRL=>AR_CTRL,BI_CTRL=>BI_CTRL,BR_CTRL=>BR_CTRL,
							OUT_MUX1=>BUS1,OUT_MUX2=>BUS2,OUT_MUX3=> BUSW);
MOLTIPLICATORE: MOL PORT MAP(CLK=>CLK,C=>C,ADD1=>BUS2,ADD2=>BUSW,RESULT=> MOL_RES_IN);
SOMMATORE: SUM PORT MAP(CLK=>CLK,A_S=>A_S,T1=>OUTMUXINVT1,T2=>OUTMUXINVT2,RESULT=>SUM_RES_IN);
REG_MOL: REG_39_M PORT MAP(CLK=>CLK,D=>MOL_RES_IN,Q=>MOL_RES_OUT);
REG_SUM : REG_40_S PORT MAP(CLK=>CLK,D=>SUM_RES_IN,Q=>SUM_RES_OUT);
R_ROUNDING: REG_ROUND PORT MAP (CLK=>CLK,ENABLE=>EN_REGR,D=>SUM_RES_OUT,Q=>REG_ROUND_OUT);
R_A1R: REG_A1R PORT MAP(CLK=>CLK,ENABLE=>EN_REGO,D=>ROUNDED(19 DOWNTO 0),Q=>A1R);
R_A1I: REG_A1I PORT MAP(CLK=>CLK,ENABLE=>EN_REGO,D=>ROUNDED(19 DOWNTO 0),Q=>A1I);
R_B1R: REG_B1R PORT MAP(CLK=>CLK,ENABLE=>EN_REGO,D=>ROUNDED(19 DOWNTO 0),Q=>B1R);
R_B1I: REG_B1I PORT MAP(CLK=>CLK,ENABLE=>EN_REGO,D=>ROUNDED(19 DOWNTO 0),Q=>B1I);
INVT1: MUX_INV PORT MAP(SEL=>SEL_INV,A=>MUXSUM_OUT,B=>MOL_RES_OUT,OUTPUT=>OUTMUXINVT1);
INVT2: MUX_INV PORT MAP(SEL=>SEL_INV,A=>MOL_RES_OUT,B=>MUXSUM_OUT,OUTPUT=>OUTMUXINVT2);

end behav;