LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all; 

ENTITY R_STONE_1 IS

PORT(
      OUTPUT_P,OUTPUT_N: OUT SIGNED(19 DOWNTO 0));
END R_STONE_1;


ARCHITECTURE BEHAV OF R_STONE_1 IS 
SIGNAL VALORE :SIGNED (19 DOWNTO 0);
BEGIN 
VALORE<= "01111111111111111111";
OUTPUT_P<=VALORE;
OUTPUT_N<= NOT VALORE;
END BEHAV;