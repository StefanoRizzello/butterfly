LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all; 

ENTITY GUARD IS

PORT ( C0AR,C1AR,C2AR,C3AR,C4AR,C5AR,C6AR,C7AR: IN SIGNED(19 downto 0);
		 C0AI,C1AI,C2AI,C3AI,C4AI,C5AI,C6AI,C7AI: IN SIGNED(19 downto 0);
		 C0BR,C1BR,C2BR,C3BR,C4BR,C5BR,C6BR,C7BR: IN SIGNED(19 downto 0);
		 C0BI,C1BI,C2BI,C3BI,C4BI,C5BI,C6BI,C7BI: IN SIGNED(19 downto 0);
		
	    C0AR_GUARD,C1AR_GUARD,C2AR_GUARD,C3AR_GUARD,C4AR_GUARD,C5AR_GUARD,C6AR_GUARD,C7AR_GUARD: 
		 OUT SIGNED(19 downto 0);
		 C0AI_GUARD,C1AI_GUARD,C2AI_GUARD,C3AI_GUARD,C4AI_GUARD,C5AI_GUARD,C6AI_GUARD,C7AI_GUARD: 
		 OUT SIGNED(19 downto 0);
		 C0BR_GUARD,C1BR_GUARD,C2BR_GUARD,C3BR_GUARD,C4BR_GUARD,C5BR_GUARD,C6BR_GUARD,C7BR_GUARD: 
		 OUT SIGNED(19 downto 0);
		 C0BI_GUARD,C1BI_GUARD,C2BI_GUARD,C3BI_GUARD,C4BI_GUARD,C5BI_GUARD,C6BI_GUARD,C7BI_GUARD: 
		 OUT SIGNED(19 downto 0));
END GUARD;

ARCHITECTURE behav OF GUARD IS

BEGIN

C0AR_GUARD(19) <= C0AR(19); C0AR_GUARD(18 DOWNTO 0) <= C0AR(19 DOWNTO 1);
C1AR_GUARD(19) <= C1AR(19); C1AR_GUARD(18 DOWNTO 0) <= C1AR(19 DOWNTO 1);
C2AR_GUARD(19) <= C2AR(19); C2AR_GUARD(18 DOWNTO 0) <= C2AR(19 DOWNTO 1);
C3AR_GUARD(19) <= C3AR(19); C3AR_GUARD(18 DOWNTO 0) <= C3AR(19 DOWNTO 1);
C4AR_GUARD(19) <= C4AR(19); C4AR_GUARD(18 DOWNTO 0) <= C4AR(19 DOWNTO 1);
C5AR_GUARD(19) <= C5AR(19); C5AR_GUARD(18 DOWNTO 0) <= C5AR(19 DOWNTO 1);
C6AR_GUARD(19) <= C6AR(19); C6AR_GUARD(18 DOWNTO 0) <= C6AR(19 DOWNTO 1);
C7AR_GUARD(19) <= C7AR(19); C7AR_GUARD(18 DOWNTO 0) <= C7AR(19 DOWNTO 1);

C0AI_GUARD(19) <= C0AI(19); C0AI_GUARD(18 DOWNTO 0) <= C0AI(19 DOWNTO 1);
C1AI_GUARD(19) <= C1AI(19); C1AI_GUARD(18 DOWNTO 0) <= C1AI(19 DOWNTO 1);
C2AI_GUARD(19) <= C2AI(19); C2AI_GUARD(18 DOWNTO 0) <= C2AI(19 DOWNTO 1);
C3AI_GUARD(19) <= C3AI(19); C3AI_GUARD(18 DOWNTO 0) <= C3AI(19 DOWNTO 1);
C4AI_GUARD(19) <= C4AI(19); C4AI_GUARD(18 DOWNTO 0) <= C4AI(19 DOWNTO 1);
C5AI_GUARD(19) <= C5AI(19); C5AI_GUARD(18 DOWNTO 0) <= C5AI(19 DOWNTO 1);
C6AI_GUARD(19) <= C6AI(19); C6AI_GUARD(18 DOWNTO 0) <= C6AI(19 DOWNTO 1);
C7AI_GUARD(19) <= C7AI(19); C7AI_GUARD(18 DOWNTO 0) <= C7AI(19 DOWNTO 1);

C0BR_GUARD(19) <= C0BR(19); C0BR_GUARD(18 DOWNTO 0) <= C0BR(19 DOWNTO 1);
C1BR_GUARD(19) <= C1BR(19); C1BR_GUARD(18 DOWNTO 0) <= C1BR(19 DOWNTO 1);
C2BR_GUARD(19) <= C2BR(19); C2BR_GUARD(18 DOWNTO 0) <= C2BR(19 DOWNTO 1);
C3BR_GUARD(19) <= C3BR(19); C3BR_GUARD(18 DOWNTO 0) <= C3BR(19 DOWNTO 1);
C4BR_GUARD(19) <= C4BR(19); C4BR_GUARD(18 DOWNTO 0) <= C4BR(19 DOWNTO 1);
C5BR_GUARD(19) <= C5BR(19); C5BR_GUARD(18 DOWNTO 0) <= C5BR(19 DOWNTO 1);
C6BR_GUARD(19) <= C6BR(19); C6BR_GUARD(18 DOWNTO 0) <= C6BR(19 DOWNTO 1);
C7BR_GUARD(19) <= C7BR(19); C7BR_GUARD(18 DOWNTO 0) <= C7BR(19 DOWNTO 1);

C0BI_GUARD(19) <= C0BI(19); C0BI_GUARD(18 DOWNTO 0) <= C0BI(19 DOWNTO 1);
C1BI_GUARD(19) <= C1BI(19); C1BI_GUARD(18 DOWNTO 0) <= C1BI(19 DOWNTO 1);
C2BI_GUARD(19) <= C2BI(19); C2BI_GUARD(18 DOWNTO 0) <= C2BI(19 DOWNTO 1);
C3BI_GUARD(19) <= C3BI(19); C3BI_GUARD(18 DOWNTO 0) <= C3BI(19 DOWNTO 1);
C4BI_GUARD(19) <= C4BI(19); C4BI_GUARD(18 DOWNTO 0) <= C4BI(19 DOWNTO 1);
C5BI_GUARD(19) <= C5BI(19); C5BI_GUARD(18 DOWNTO 0) <= C5BI(19 DOWNTO 1);
C6BI_GUARD(19) <= C6BI(19); C6BI_GUARD(18 DOWNTO 0) <= C6BI(19 DOWNTO 1);
C7BI_GUARD(19) <= C7BI(19); C7BI_GUARD(18 DOWNTO 0) <= C7BI(19 DOWNTO 1);



END behav;