LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all; 

ENTITY REG_SEQ IS

PORT (CLK,D0,D1,D2,D3,SET,RESET,EN0,EN1,EN2,EN3: IN STD_LOGIC;
		Q0,Q1,Q2,Q3: OUT STD_LOGIC);		 
END REG_SEQ;

ARCHITECTURE behav OF REG_SEQ IS

COMPONENT FF_SEQ IS
PORT (CLK,D,SET,RESET,ENABLE: IN STD_LOGIC;
		Q: OUT STD_LOGIC);		 
END COMPONENT;


BEGIN

FF0: FF_SEQ PORT MAP(CLK=>CLK,D=>D0,SET=>SET,RESET=>RESET,ENABLE=>EN0,Q=>Q0);
FF1: FF_SEQ PORT MAP(CLK=>CLK,D=>D1,SET=>SET,RESET=>RESET,ENABLE=>EN1,Q=>Q1);
FF2: FF_SEQ PORT MAP(CLK=>CLK,D=>D2,SET=>SET,RESET=>RESET,ENABLE=>EN2,Q=>Q2);
FF3: FF_SEQ PORT MAP(CLK=>CLK,D=>D3,SET=>SET,RESET=>RESET,ENABLE=>EN3,Q=>Q3);


END behav;