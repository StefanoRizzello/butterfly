LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all; 

ENTITY FFT_16 IS

PORT ( CLK,RESET: IN STD_LOGIC;
		 DONE,READY: OUT STD_LOGIC;
       C0AR,C1AR,C2AR,C3AR,C4AR,C5AR,C6AR,C7AR: IN SIGNED(19 downto 0);
		 C0AI,C1AI,C2AI,C3AI,C4AI,C5AI,C6AI,C7AI: IN SIGNED(19 downto 0);
		 C0BR,C1BR,C2BR,C3BR,C4BR,C5BR,C6BR,C7BR: IN SIGNED(19 downto 0);
		 C0BI,C1BI,C2BI,C3BI,C4BI,C5BI,C6BI,C7BI: IN SIGNED(19 downto 0);
		
	    C0AR_OUT,C1AR_OUT,C2AR_OUT,C3AR_OUT,C4AR_OUT,C5AR_OUT,C6AR_OUT,C7AR_OUT: 
		 OUT SIGNED(19 downto 0);
		 C0AI_OUT,C1AI_OUT,C2AI_OUT,C3AI_OUT,C4AI_OUT,C5AI_OUT,C6AI_OUT,C7AI_OUT: 
		 OUT SIGNED(19 downto 0);
		 C0BR_OUT,C1BR_OUT,C2BR_OUT,C3BR_OUT,C4BR_OUT,C5BR_OUT,C6BR_OUT,C7BR_OUT: 
		 OUT SIGNED(19 downto 0);
		 C0BI_OUT,C1BI_OUT,C2BI_OUT,C3BI_OUT,C4BI_OUT,C5BI_OUT,C6BI_OUT,C7BI_OUT: 
		 OUT SIGNED(19 downto 0));
       
		 
END FFT_16;

ARCHITECTURE behav OF FFT_16 IS

COMPONENT BF IS
PORT ( CLK, ENABLE: IN std_logic;
       AI,AR,BI,BR,WR,WI: IN SIGNED(19 downto 0); -- va cambiato il formato e conversioni
      SEL_INV,SEL3,SEL1,SELSUM,C,A_S,EN_REGR : IN std_logic;
		SEL2: IN std_logic_vector(1 downto 0);
		EN_REGO: IN std_logic_vector(2 downto 0);
		A1R,A1I,B1R,B1I,AI_CTRL,AR_CTRL,BI_CTRL,BR_CTRL: OUT SIGNED(19 downto 0));
END COMPONENT;

COMPONENT OR_PORT IS
PORT ( B0AR,B1AR,B2AR,B3AR,B4AR,B5AR,B6AR,B7AR: IN SIGNED(19 downto 0);
		 B0AI,B1AI,B2AI,B3AI,B4AI,B5AI,B6AI,B7AI: IN SIGNED(19 downto 0);
		 B0BR,B1BR,B2BR,B3BR,B4BR,B5BR,B6BR,B7BR: IN SIGNED(19 downto 0);
		 B0BI,B1BI,B2BI,B3BI,B4BI,B5BI,B6BI,B7BI: IN SIGNED(19 downto 0);
       START: OUT std_logic);
END COMPONENT;

COMPONENT XOR_CHECK IS
PORT ( B0AR,B1AR,B2AR,B3AR,B4AR,B5AR,B6AR,B7AR: IN SIGNED(19 downto 0);
		 B0AI,B1AI,B2AI,B3AI,B4AI,B5AI,B6AI,B7AI: IN SIGNED(19 downto 0);
		 B0BR,B1BR,B2BR,B3BR,B4BR,B5BR,B6BR,B7BR: IN SIGNED(19 downto 0);
		 B0BI,B1BI,B2BI,B3BI,B4BI,B5BI,B6BI,B7BI: IN SIGNED(19 downto 0);
		
	    B0AR_OLD,B1AR_OLD,B2AR_OLD,B3AR_OLD,B4AR_OLD,B5AR_OLD,B6AR_OLD,B7AR_OLD: 
		 IN SIGNED(19 downto 0);
		 B0AI_OLD,B1AI_OLD,B2AI_OLD,B3AI_OLD,B4AI_OLD,B5AI_OLD,B6AI_OLD,B7AI_OLD: 
		 IN SIGNED(19 downto 0);
		 B0BR_OLD,B1BR_OLD,B2BR_OLD,B3BR_OLD,B4BR_OLD,B5BR_OLD,B6BR_OLD,B7BR_OLD: 
		 IN SIGNED(19 downto 0);
		 B0BI_OLD,B1BI_OLD,B2BI_OLD,B3BI_OLD,B4BI_OLD,B5BI_OLD,B6BI_OLD,B7BI_OLD: 
		 IN SIGNED(19 downto 0);
       
		 OUT_XOR_CHECK: OUT std_logic);
END COMPONENT;	

COMPONENT R_STONE_0 IS
PORT(
      OUTPUT: OUT SIGNED(19 DOWNTO 0));
END COMPONENT;	 

COMPONENT R_STONE_1 IS
PORT(
      OUTPUT_P,OUTPUT_N: OUT SIGNED(19 DOWNTO 0));
END COMPONENT;

COMPONENT R_STONE_3 IS
PORT(
      OUTPUT_P,OUTPUT_N: OUT SIGNED(19 DOWNTO 0));
END COMPONENT;

COMPONENT R_STONE_7 IS
PORT(
      OUTPUT_P,OUTPUT_N: OUT SIGNED(19 DOWNTO 0));
END COMPONENT;

COMPONENT R_STONE_9 IS
PORT(
      OUTPUT_P,OUTPUT_N: OUT SIGNED(19 DOWNTO 0));
END COMPONENT;

COMPONENT CU_BF IS
PORT( LOAD,SEQ,CLK,RESET: IN std_logic;
		CTRL_OUT: OUT std_logic_vector(14 downto 0));
END COMPONENT;

COMPONENT CU_TOP IS 
PORT( START,PROGRESS,FREE_M,END_BF,SEQ,CLK,RESET: IN std_logic;
		CTRL_TOP_OUT: OUT std_logic_vector(5 downto 0));
END COMPONENT;

COMPONENT start_sense IS 
PORT (D, CLK,set,enable : IN std_logic;
       SENSE : OUT std_logic);
END  COMPONENT;

COMPONENT REG_STATUS IS 
PORT ( CLK,set,enable0,enable1,enable2,enable3,RESET : IN std_logic;
       Q_OUT: OUT std_logic_vector (3 downto 0));
END  COMPONENT;

COMPONENT REG_SEQ IS
PORT (CLK,D0,D1,D2,D3,SET,RESET,EN0,EN1,EN2,EN3: IN STD_LOGIC;
		Q0,Q1,Q2,Q3: OUT STD_LOGIC);		 
END COMPONENT;
		
COMPONENT GUARD IS
PORT ( C0AR,C1AR,C2AR,C3AR,C4AR,C5AR,C6AR,C7AR: IN SIGNED(19 downto 0);
		 C0AI,C1AI,C2AI,C3AI,C4AI,C5AI,C6AI,C7AI: IN SIGNED(19 downto 0);
		 C0BR,C1BR,C2BR,C3BR,C4BR,C5BR,C6BR,C7BR: IN SIGNED(19 downto 0);
		 C0BI,C1BI,C2BI,C3BI,C4BI,C5BI,C6BI,C7BI: IN SIGNED(19 downto 0);
		
	    C0AR_GUARD,C1AR_GUARD,C2AR_GUARD,C3AR_GUARD,C4AR_GUARD,C5AR_GUARD,C6AR_GUARD,C7AR_GUARD: 
		 OUT SIGNED(19 downto 0);
		 C0AI_GUARD,C1AI_GUARD,C2AI_GUARD,C3AI_GUARD,C4AI_GUARD,C5AI_GUARD,C6AI_GUARD,C7AI_GUARD: 
		 OUT SIGNED(19 downto 0);
		 C0BR_GUARD,C1BR_GUARD,C2BR_GUARD,C3BR_GUARD,C4BR_GUARD,C5BR_GUARD,C6BR_GUARD,C7BR_GUARD: 
		 OUT SIGNED(19 downto 0);
		 C0BI_GUARD,C1BI_GUARD,C2BI_GUARD,C3BI_GUARD,C4BI_GUARD,C5BI_GUARD,C6BI_GUARD,C7BI_GUARD: 
		 OUT SIGNED(19 downto 0));
END COMPONENT;	
		
-- SEGNALI CTRL TOP OUT
SIGNAL FF_VALUE_S,EN_FF_S: STD_LOGIC;
SIGNAL RESET_OUT: STD_LOGIC;
SIGNAL PROGRESS_S: STD_LOGIC_VECTOR (3 downto 0);

SIGNAL EN_REGS0,EN_REGS1,EN_REGS2,EN_REGS3,FREE_M_S: STD_LOGIC;

SIGNAL NEW_PROGRESS_S : STD_LOGIC;


-- SEGNALI PER LA CU DELLE BF USCITA
SIGNAL SEL3_S0,SEL1_S0,SELSUM_S0,C_S0,A_S_S0,EN_REGR_S0,ENABLE_S0,SEL_INV_S0 : STD_LOGIC; 
SIGNAL SEL3_S1,SEL1_S1,SELSUM_S1,C_S1,A_S_S1,EN_REGR_S1,ENABLE_S1,SEL_INV_S1 : STD_LOGIC;
SIGNAL SEL3_S2,SEL1_S2,SELSUM_S2,C_S2,A_S_S2,EN_REGR_S2,ENABLE_S2,SEL_INV_S2 : STD_LOGIC;
SIGNAL SEL3_S3,SEL1_S3,SELSUM_S3,C_S3,A_S_S3,EN_REGR_S3,ENABLE_S3,SEL_INV_S3 : STD_LOGIC;

SIGNAL SEL2_S0: STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL SEL2_S1: STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL SEL2_S2: STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL SEL2_S3: STD_LOGIC_VECTOR(1 DOWNTO 0);

SIGNAL EN_REGO_S0: STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL EN_REGO_S1: STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL EN_REGO_S2: STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL EN_REGO_S3: STD_LOGIC_VECTOR(2 DOWNTO 0);

--SEGNALI PER LA CU TOP INGRESSO
SIGNAL START_S,START_S_TOP, OUT_XOR_CHECK_S,NEW_OUT_XOR_CHECK_S : STD_LOGIC;
SIGNAL END_BF_TOP,FREE_M_TOP : STD_LOGIC;

-- SONO I SEGNALI DA MANDARE AI REGISTRI WR WI
SIGNAL  P_0,P_1,P_3,P_7,P_9 : SIGNED (19 DOWNTO 0); 
SIGNAL  N_1,N_3,N_7,N_9 :SIGNED (19 DOWNTO 0);

-- SEGNALI PER CONTROLLO XOR (da mettere tra step 0 e XOR_CHECK
SIGNAL AI0_CTRL,AI1_CTRL,AI2_CTRL,AI3_CTRL,AI4_CTRL,AI5_CTRL,AI6_CTRL,AI7_CTRL : SIGNED (19 DOWNTO 0);
SIGNAL AR0_CTRL,AR1_CTRL,AR2_CTRL,AR3_CTRL,AR4_CTRL,AR5_CTRL,AR6_CTRL,AR7_CTRL : SIGNED (19 DOWNTO 0);
SIGNAL BR0_CTRL,BR1_CTRL,BR2_CTRL,BR3_CTRL,BR4_CTRL,BR5_CTRL,BR6_CTRL,BR7_CTRL : SIGNED (19 DOWNTO 0);
SIGNAL BI0_CTRL,BI1_CTRL,BI2_CTRL,BI3_CTRL,BI4_CTRL,BI5_CTRL,BI6_CTRL,BI7_CTRL : SIGNED (19 DOWNTO 0);

-- SEGNALI PER COLLEGARE UNA BF ALLA SUCCESSIVA
SIGNAL S01_0_AR,S01_1_AR, S01_2_AR, S01_3_AR, S01_4_AR, S01_5_AR, S01_6_AR, S01_7_AR:SIGNED(19 DOWNTO 0);
SIGNAL S01_0_AI,S01_1_AI, S01_2_AI, S01_3_AI, S01_4_AI, S01_5_AI, S01_6_AI, S01_7_AI:SIGNED(19 DOWNTO 0);
SIGNAL S01_0_BR,S01_1_BR, S01_2_BR, S01_3_BR, S01_4_BR, S01_5_BR, S01_6_BR, S01_7_BR:SIGNED(19 DOWNTO 0); 
SIGNAL S01_0_BI,S01_1_BI, S01_2_BI, S01_3_BI, S01_4_BI, S01_5_BI, S01_6_BI, S01_7_BI:SIGNED(19 DOWNTO 0);

SIGNAL S12_0_AR,S12_1_AR, S12_2_AR, S12_3_AR, S12_4_AR, S12_5_AR, S12_6_AR, S12_7_AR:SIGNED(19 DOWNTO 0);
SIGNAL S12_0_AI,S12_1_AI, S12_2_AI, S12_3_AI, S12_4_AI, S12_5_AI, S12_6_AI, S12_7_AI:SIGNED(19 DOWNTO 0);
SIGNAL S12_0_BR,S12_1_BR, S12_2_BR, S12_3_BR, S12_4_BR, S12_5_BR, S12_6_BR, S12_7_BR:SIGNED(19 DOWNTO 0); 
SIGNAL S12_0_BI,S12_1_BI, S12_2_BI, S12_3_BI, S12_4_BI, S12_5_BI, S12_6_BI, S12_7_BI:SIGNED(19 DOWNTO 0);

SIGNAL S23_0_AR,S23_1_AR, S23_2_AR, S23_3_AR, S23_4_AR, S23_5_AR, S23_6_AR, S23_7_AR:SIGNED(19 DOWNTO 0);
SIGNAL S23_0_AI,S23_1_AI, S23_2_AI, S23_3_AI, S23_4_AI, S23_5_AI, S23_6_AI, S23_7_AI:SIGNED(19 DOWNTO 0);
SIGNAL S23_0_BR,S23_1_BR, S23_2_BR, S23_3_BR, S23_4_BR, S23_5_BR, S23_6_BR, S23_7_BR:SIGNED(19 DOWNTO 0);
SIGNAL S23_0_BI,S23_1_BI, S23_2_BI, S23_3_BI, S23_4_BI, S23_5_BI, S23_6_BI, S23_7_BI:SIGNED(19 DOWNTO 0);

-- GUARD BIT
SIGNAL C0AR_GUARD_S,C1AR_GUARD_S,C2AR_GUARD_S,C3AR_GUARD_S,C4AR_GUARD_S,C5AR_GUARD_S,C6AR_GUARD_S,C7AR_GUARD_S : SIGNED(19 DOWNTO 0);
SIGNAL C0AI_GUARD_S,C1AI_GUARD_S,C2AI_GUARD_S,C3AI_GUARD_S,C4AI_GUARD_S,C5AI_GUARD_S,C6AI_GUARD_S,C7AI_GUARD_S : SIGNED(19 DOWNTO 0);
SIGNAL C0BR_GUARD_S,C1BR_GUARD_S,C2BR_GUARD_S,C3BR_GUARD_S,C4BR_GUARD_S,C5BR_GUARD_S,C6BR_GUARD_S,C7BR_GUARD_S : SIGNED(19 DOWNTO 0);
SIGNAL C0BI_GUARD_S,C1BI_GUARD_S,C2BI_GUARD_S,C3BI_GUARD_S,C4BI_GUARD_S,C5BI_GUARD_S,C6BI_GUARD_S,C7BI_GUARD_S : SIGNED(19 DOWNTO 0);


SIGNAL SENSE_S: STD_LOGIC;

SIGNAL SEQ_CU0,SEQ_CU1,SEQ_CU2,SEQ_CU3: STD_LOGIC;

SIGNAL SET_FALSO: STD_LOGIC;

SIGNAL SET_REG_SEQ: STD_LOGIC;

BEGIN 


SET_REG_SEQ <= FF_VALUE_S AND NEW_OUT_XOR_CHECK_S;
NEW_OUT_XOR_CHECK_S <= OUT_XOR_CHECK_S AND START_S;
SET_FALSO <= RESET_OUT AND FF_VALUE_S; 
START_S_TOP <= SENSE_S AND START_S;
NEW_PROGRESS_S <= PROGRESS_S(3) OR PROGRESS_S(2) OR PROGRESS_S(1) OR PROGRESS_S(0);

-- BF DELLO STEP 0 COLLEGATE DIRETTAMENTI AGLI INGRESSI DELLA FFT 16
BF_0_0: BF PORT MAP(AI=>C0AI_GUARD_S,AR=>C0AR_GUARD_S,BR=>C0BR_GUARD_S,BI=>C0BI_GUARD_S, A1R=>S01_0_AR,A1I=>S01_0_AI,B1R=>S01_0_BR,B1I=>							S01_0_BI,SEL3=> SEL3_S0,SEL1=>SEL1_S0,SELSUM=>SELSUM_S0,C=>C_S0,A_S=>A_S_S0,EN_REGR=>							EN_REGR_S0,ENABLE=>ENABLE_S0,SEL2=> SEL2_S0,EN_REGO=>EN_REGO_S0,WR=>P_1,WI=>P_0,CLK=>CLK,AI_CTRL=>AI1_CTRL,AR_CTRL=>AR0_CTRL,BI_CTRL=>BI0_CTRL,BR_CTRL=>BR0_CTRL,SEL_INV=>SEL_INV_S0);
BF_0_1: BF PORT MAP(AI=>C1AI_GUARD_S,AR=>C1AR_GUARD_S,BR=>C1BR_GUARD_S,BI=>C1BI_GUARD_S, A1R=>S01_1_AR,A1I=>S01_1_AI,B1R=>S01_1_BR,B1I=>							S01_1_BI, SEL3=> SEL3_S0,SEL1=>SEL1_S0,SELSUM=>SELSUM_S0,C=>C_S0,A_S=>A_S_S0,EN_REGR=>							EN_REGR_S0,ENABLE=>ENABLE_S0,SEL2=> SEL2_S0,EN_REGO=>EN_REGO_S0,WR=>P_1,WI=>P_0, CLK=>CLK,AI_CTRL=>AI0_CTRL,AR_CTRL=>AR1_CTRL,BI_CTRL=>BI1_CTRL,BR_CTRL=>BR1_CTRL,SEL_INV=>SEL_INV_S0);
BF_0_2: BF PORT MAP(AI=>C2AI_GUARD_S,AR=>C2AR_GUARD_S,BR=>C2BR_GUARD_S,BI=>C2BI_GUARD_S, A1R=>S01_2_AR,A1I=>S01_2_AI,B1R=>S01_2_BR,B1I=>							S01_2_BI,SEL3=> SEL3_S0,SEL1=>SEL1_S0,SELSUM=>SELSUM_S0,C=>C_S0,A_S=>A_S_S0,							EN_REGR=>EN_REGR_S0,ENABLE=>ENABLE_S0,SEL2=> SEL2_S0,EN_REGO=>EN_REGO_S0,WR=>P_1,WI=>P_0,CLK=>CLK,AI_CTRL=>AI2_CTRL,AR_CTRL=>AR2_CTRL,BI_CTRL=>BI2_CTRL,BR_CTRL=>BR2_CTRL,SEL_INV=>SEL_INV_S0);
BF_0_3: BF PORT MAP(AI=>C3AI_GUARD_S,AR=>C3AR_GUARD_S,BR=>C3BR_GUARD_S,BI=>C3BI_GUARD_S, A1R=>S01_3_AR,A1I=>S01_3_AI,B1R=>S01_3_BR,B1I=>							S01_3_BI,SEL3=> SEL3_S0,SEL1=>SEL1_S0,SELSUM=>SELSUM_S0,C=>C_S0,A_S=>A_S_S0,EN_REGR=>							EN_REGR_S0,ENABLE=>ENABLE_S0,SEL2=> SEL2_S0,EN_REGO=>EN_REGO_S0,WR=>P_1,WI=>P_0, CLK=>CLK,AI_CTRL=>AI3_CTRL,AR_CTRL=>AR3_CTRL,BI_CTRL=>BI3_CTRL,BR_CTRL=>BR3_CTRL,SEL_INV=>SEL_INV_S0);
BF_0_4: BF PORT MAP(AI=>C4AI_GUARD_S,AR=>C4AR_GUARD_S,BR=>C4BR_GUARD_S,BI=>C4BI_GUARD_S, A1R=>S01_4_AR,A1I=>S01_4_AI,B1R=>S01_4_BR,B1I=>							S01_4_BI, SEL3=> SEL3_S0,SEL1=>SEL1_S0,SELSUM=>SELSUM_S0,C=>C_S0,A_S=>A_S_S0,EN_REGR=>							EN_REGR_S0,ENABLE=>ENABLE_S0,SEL2=> SEL2_S0,EN_REGO=>EN_REGO_S0,WR=>P_1,WI=>P_0, CLK=>CLK,AI_CTRL=>AI4_CTRL,AR_CTRL=>AR4_CTRL,BI_CTRL=>BI4_CTRL,BR_CTRL=>BR4_CTRL,SEL_INV=>SEL_INV_S0);
BF_0_5: BF PORT MAP(AI=>C5AI_GUARD_S,AR=>C5AR_GUARD_S,BR=>C5BR_GUARD_S,BI=>C5BI_GUARD_S, A1R=>S01_5_AR,A1I=>S01_5_AI,B1R=>S01_5_BR,B1I=>							S01_5_BI, SEL3=> SEL3_S0,SEL1=>SEL1_S0,SELSUM=>SELSUM_S0,C=>C_S0,A_S=>A_S_S0,							EN_REGR=>EN_REGR_S0,ENABLE=>ENABLE_S0,SEL2=> SEL2_S0,EN_REGO=>EN_REGO_S0,WR=>P_1,WI=>P_0,CLK=>CLK,AI_CTRL=>AI5_CTRL,AR_CTRL=>AR5_CTRL,BI_CTRL=>BI5_CTRL,BR_CTRL=>BR5_CTRL,SEL_INV=>SEL_INV_S0);
BF_0_6: BF PORT MAP(AI=>C6AI_GUARD_S,AR=>C6AR_GUARD_S,BR=>C6BR_GUARD_S,BI=>C6BI_GUARD_S, A1R=>S01_6_AR,A1I=>S01_6_AI,B1R=>S01_6_BR,B1I=>							S01_6_BI, SEL3=> SEL3_S0,SEL1=>SEL1_S0,SELSUM=>SELSUM_S0,C=>C_S0,A_S=>A_S_S0,EN_REGR=>							EN_REGR_S0,ENABLE=>ENABLE_S0,SEL2=> SEL2_S0,EN_REGO=>EN_REGO_S0,WR=>P_1,WI=>P_0, CLK=>CLK,AI_CTRL=>AI6_CTRL,AR_CTRL=>AR6_CTRL,BI_CTRL=>BI6_CTRL,BR_CTRL=>BR6_CTRL,SEL_INV=>SEL_INV_S0);
BF_0_7: BF PORT MAP(AI=>C7AI_GUARD_S,AR=>C7AR_GUARD_S,BR=>C7BR_GUARD_S,BI=>C7BI_GUARD_S, A1R=>S01_7_AR,A1I=>S01_7_AI,B1R=>S01_7_BR,B1I=>							S01_7_BI, SEL3=> SEL3_S0,SEL1=>SEL1_S0,SELSUM=>SELSUM_S0,C=>C_S0,A_S=>A_S_S0,EN_REGR=>							EN_REGR_S0,ENABLE=>ENABLE_S0,SEL2=> SEL2_S0,EN_REGO=>EN_REGO_S0,WR=>P_1,WI=>P_0, CLK=>CLK,AI_CTRL=>AI7_CTRL,AR_CTRL=>AR7_CTRL,BI_CTRL=>BI7_CTRL,BR_CTRL=>BR7_CTRL,SEL_INV=>SEL_INV_S0);

-- BF STEP 1

BF_1_0: BF PORT MAP(AI=>S01_0_AI,AR=>S01_0_AR,BR=>S01_4_AR,BI=>S01_4_AI, A1R=>S12_0_AR,A1I=>S12_0_AI,B1R=>							S12_0_BR,B1I=>S12_0_BI,SEL3=>SEL3_S1,SEL1=>SEL1_S1,SELSUM=>SELSUM_S1,C=>C_S1,A_S=>							A_S_S1,EN_REGR=>EN_REGR_S1,ENABLE=>ENABLE_S1,SEL2=> SEL2_S1,EN_REGO=>EN_REGO_S1,WR=>P_1,WI=>P_0, CLK=>CLK,SEL_INV=>SEL_INV_S1);
BF_1_1: BF PORT MAP(AI=>S01_1_AI,AR=>S01_1_AR,BR=>S01_5_AR,BI=>S01_5_AI, A1R=>S12_1_AR,A1I=>S12_1_AI,B1R=>							S12_1_BR,B1I=>S12_1_BI,SEL3=>SEL3_S1,SEL1=>	SEL1_S1,SELSUM=>SELSUM_S1,C=>C_S1,A_S							=>	A_S_S1,EN_REGR=>EN_REGR_S1,ENABLE=>ENABLE_S1,SEL2=> SEL2_S1,EN_REGO=>EN_REGO_S1,WR=>P_1,WI=>P_0, CLK=>CLK,SEL_INV=>SEL_INV_S1);
BF_1_2: BF PORT MAP(AI=>S01_2_AI,AR=>S01_2_AR,BR=>S01_6_AR,BI=>S01_6_AI, A1R=>S12_2_AR,A1I=>S12_2_AI,B1R=>							S12_2_BR,B1I=>S12_2_BI,SEL3=>SEL3_S1,SEL1=>SEL1_S1,SELSUM=>SELSUM_S1,C=>C_S1,A_S=>							A_S_S1,EN_REGR=>EN_REGR_S1,ENABLE=>ENABLE_S1,SEL2=> SEL2_S1,EN_REGO=>EN_REGO_S1,WR=>P_1,WI=>P_0, CLK=>CLK,SEL_INV=>SEL_INV_S1);
BF_1_3: BF PORT MAP(AI=>S01_3_AI,AR=>S01_3_AR,BR=>S01_7_AR,BI=>S01_7_AI, A1R=>S12_3_AR,A1I=>S12_3_AI,B1R=>							S12_3_BR,B1I=>S12_3_BI,SEL3=>SEL3_S1,SEL1=>SEL1_S1,SELSUM=>SELSUM_S1,C=>C_S1,A_S=>							A_S_S1,EN_REGR=>EN_REGR_S1,ENABLE=>ENABLE_S1,SEL2=> SEL2_S1,EN_REGO=>EN_REGO_S1,WR=>P_1,WI=>P_0, CLK=>CLK,SEL_INV=>SEL_INV_S1);
BF_1_4: BF PORT MAP(AI=>S01_0_BI,AR=>S01_0_BR,BR=>S01_4_BR,BI=>S01_4_BI, A1R=>S12_4_AR,A1I=>S12_4_AI,B1R=>							S12_4_BR,B1I=>S12_4_BI,SEL3=>SEL3_S1,SEL1=>	SEL1_S1,SELSUM=>SELSUM_S1,C=>C_S1,A_S=>							A_S_S1,EN_REGR=>EN_REGR_S1,ENABLE=>ENABLE_S1,SEL2=> SEL2_S1,EN_REGO=>EN_REGO_S1,WR=>P_0,WI=>N_1, CLK=>CLK,SEL_INV=>SEL_INV_S1);
BF_1_5: BF PORT MAP(AI=>S01_1_BI,AR=>S01_1_BR,BR=>S01_5_BR,BI=>S01_5_BI, A1R=>S12_5_AR,A1I=>S12_5_AI,B1R=>							S12_5_BR,B1I=>S12_5_BI,SEL3=>SEL3_S1,SEL1=>SEL1_S1,SELSUM=>SELSUM_S1,C=>C_S1,A_S=>							A_S_S1,EN_REGR=>EN_REGR_S1,ENABLE=>ENABLE_S1,SEL2=> SEL2_S1,EN_REGO=>EN_REGO_S1,WR=>P_0,WI=>N_1, CLK=>CLK,SEL_INV=>SEL_INV_S1);
BF_1_6: BF PORT MAP(AI=>S01_2_BI,AR=>S01_2_BR,BR=>S01_6_BR,BI=>S01_6_BI, A1R=>S12_6_AR,A1I=>S12_6_AI,B1R=>							S12_6_BR,B1I=>S12_6_BI,SEL3=>SEL3_S1,SEL1=>SEL1_S1,SELSUM=>SELSUM_S1,C=>C_S1,A_S=>							A_S_S1,EN_REGR=>EN_REGR_S1,ENABLE=>ENABLE_S1,SEL2=> SEL2_S1,EN_REGO=>EN_REGO_S1,WR=>P_0,WI=>N_1, CLK=>CLK,SEL_INV=>SEL_INV_S1);
BF_1_7: BF PORT MAP(AI=>S01_3_BI,AR=>S01_3_BR,BR=>S01_7_BR,BI=>S01_7_BI, A1R=>S12_7_AR,A1I=>S12_7_AI,B1R=>							S12_7_BR,B1I=>S12_7_BI,SEL3=>SEL3_S1,SEL1=>SEL1_S1,SELSUM=>SELSUM_S1,C=>C_S1,A_S=>							A_S_S1,EN_REGR=>EN_REGR_S1,ENABLE=>ENABLE_S1,SEL2=> SEL2_S1,EN_REGO=>EN_REGO_S1,WR=>P_0,WI=>N_1, CLK=>CLK,SEL_INV=>SEL_INV_S1);

-- BF STEP 2

BF_2_0: BF PORT MAP(AI=>S12_0_AI,AR=>S12_0_AR,BR=>S12_2_AR,BI=>S12_2_AI, A1R=>S23_0_AR,A1I=>S23_0_AI,B1R=>							S23_0_BR,B1I=>S23_0_BI,SEL3=>SEL3_S2,SEL1=>SEL1_S2,SELSUM=>SELSUM_S2,C=>C_S2,A_S=>							A_S_S2,EN_REGR=>EN_REGR_S2,ENABLE=>ENABLE_S2,SEL2=> SEL2_S2,EN_REGO=>EN_REGO_S2,WR=>P_1,WI=>P_0, CLK=>CLK,SEL_INV=>SEL_INV_S2);
BF_2_1: BF PORT MAP(AI=>S12_1_AI,AR=>S12_1_AR,BR=>S12_3_AR,BI=>S12_3_AI, A1R=>S23_1_AR,A1I=>S23_1_AI,B1R=>							S23_1_BR,B1I=>S23_1_BI,SEL3=>SEL3_S2,SEL1=>SEL1_S2,SELSUM=>SELSUM_S2,C=>C_S2,A_S=>							A_S_S2,EN_REGR=>EN_REGR_S2,ENABLE=>ENABLE_S2,SEL2=> SEL2_S2,EN_REGO=>EN_REGO_S2,WR=>P_1,WI=>P_0, CLK=>CLK,SEL_INV=>SEL_INV_S2);
BF_2_2: BF PORT MAP(AI=>S12_0_BI,AR=>S12_0_BR,BR=>S12_2_BR,BI=>S12_2_BI, A1R=>S23_2_AR,A1I=>S23_2_AI,B1R=>							S23_2_BR,B1I=>S23_2_BI,SEL3=>SEL3_S2,SEL1=>SEL1_S2,SELSUM=>SELSUM_S2,C=>C_S2,A_S=>							A_S_S2,EN_REGR=>EN_REGR_S2,ENABLE=>ENABLE_S2,SEL2=> SEL2_S2,EN_REGO=>EN_REGO_S2,WR=>P_0,WI=>N_1, CLK=>CLK,SEL_INV=>SEL_INV_S2);
BF_2_3: BF PORT MAP(AI=>S12_1_BI,AR=>S12_1_BR,BR=>S12_3_BR,BI=>S12_3_BI, A1R=>S23_3_AR,A1I=>S23_3_AI,B1R=>							S23_3_BR,B1I=>S23_3_BI,SEL3=>SEL3_S2,SEL1=>SEL1_S2,SELSUM=>SELSUM_S2,C=>C_S2,A_S=>							A_S_S2,EN_REGR=>EN_REGR_S2,ENABLE=>ENABLE_S2,SEL2=> SEL2_S2,EN_REGO=>EN_REGO_S2,WR=>P_0,WI=>N_1, CLK=>CLK,SEL_INV=>SEL_INV_S2);
BF_2_4: BF PORT MAP(AI=>S12_4_AI,AR=>S12_4_AR,BR=>S12_6_AR,BI=>S12_6_AI, A1R=>S23_4_AR,A1I=>S23_4_AI,B1R=>							S23_4_BR,B1I=>S23_4_BI,SEL3=>SEL3_S2,SEL1=>SEL1_S2,SELSUM=>SELSUM_S2,C=>C_S2,A_S=>							A_S_S2,EN_REGR=>EN_REGR_S2,ENABLE=>ENABLE_S2,SEL2=> SEL2_S2,EN_REGO=>EN_REGO_S2,WR=>P_7,WI=>N_7, CLK=>CLK,SEL_INV=>SEL_INV_S2);
BF_2_5: BF PORT MAP(AI=>S12_5_AI,AR=>S12_5_AR,BR=>S12_7_AR,BI=>S12_7_AI, A1R=>S23_5_AR,A1I=>S23_5_AI,B1R=>							S23_5_BR,B1I=>S23_5_BI,SEL3=>SEL3_S2,SEL1=>SEL1_S2,SELSUM=>SELSUM_S2,C=>C_S2,A_S=>							A_S_S2,EN_REGR=>EN_REGR_S2,ENABLE=>ENABLE_S2,SEL2=> SEL2_S2,EN_REGO=>EN_REGO_S2,WR=>P_7,WI=>N_7, CLK=>CLK,SEL_INV=>SEL_INV_S2);
BF_2_6: BF PORT MAP(AI=>S12_4_BI,AR=>S12_4_BR,BR=>S12_6_BR,BI=>S12_6_BI, A1R=>S23_6_AR,A1I=>S23_6_AI,B1R=>							S23_6_BR,B1I=>S23_6_BI,SEL3=>SEL3_S2,SEL1=>SEL1_S2,SELSUM=>SELSUM_S2,C=>C_S2,A_S=>							A_S_S2,EN_REGR=>EN_REGR_S2,ENABLE=>ENABLE_S2,SEL2=> SEL2_S2,EN_REGO=>EN_REGO_S2,WR=>N_7,WI=>N_7, CLK=>CLK,SEL_INV=>SEL_INV_S2);
BF_2_7: BF PORT MAP(AI=>S12_5_BI,AR=>S12_5_BR,BR=>S12_7_BR,BI=>S12_7_BI, A1R=>S23_7_AR,A1I=>S23_7_AI,B1R=>							S23_7_BR,B1I=>S23_7_BI,SEL3=>SEL3_S2,SEL1=>SEL1_S2,SELSUM=>SELSUM_S2,C=>C_S2,A_S=>							A_S_S2,EN_REGR=>EN_REGR_S2,ENABLE=>ENABLE_S2,SEL2=> SEL2_S2,EN_REGO=>EN_REGO_S2,WR=>N_7,WI=>N_7, CLK=>CLK,SEL_INV=>SEL_INV_S2);

-- BF STEP 3 (ULTIMO)

BF_3_0: BF PORT MAP(AI=>S23_0_AI,AR=>S23_0_AR,BR=>S23_1_AR,BI=>S23_1_AI, A1R=>C0AR_OUT,A1I=>C0AI_OUT,B1R=>							C0BR_OUT,B1I=>C0BI_OUT,SEL3=>SEL3_S3,SEL1=>SEL1_S3,SELSUM=>SELSUM_S3,C=>C_S3,A_S=>							A_S_S3,EN_REGR=>EN_REGR_S3,ENABLE=>ENABLE_S3,SEL2=> SEL2_S3,EN_REGO=>EN_REGO_S3,WR=>P_1,WI=>P_0, CLK=>CLK,SEL_INV=>SEL_INV_S3);
BF_3_1: BF PORT MAP(AI=>S23_0_BI,AR=>S23_0_BR,BR=>S23_1_BR,BI=>S23_1_BI, A1R=>C1AR_OUT,A1I=>C1AI_OUT,B1R=>							C1BR_OUT,B1I=>C1BI_OUT,SEL3=>SEL3_S3,SEL1=>SEL1_S3,SELSUM=>SELSUM_S3,C=>C_S3,A_S=>							A_S_S3,EN_REGR=>EN_REGR_S3,ENABLE=>ENABLE_S3,SEL2=> SEL2_S3,EN_REGO=>EN_REGO_S3,WR=>P_0,WI=>N_1, CLK=>CLK,SEL_INV=>SEL_INV_S3);
BF_3_2: BF PORT MAP(AI=>S23_2_AI,AR=>S23_2_AR,BR=>S23_3_AR,BI=>S23_3_AI, A1R=>C2AR_OUT,A1I=>C2AI_OUT,B1R=>							C2BR_OUT,B1I=>C2BI_OUT,SEL3=>SEL3_S3,SEL1=>SEL1_S3,SELSUM=>SELSUM_S3,C=>C_S3,A_S=>							A_S_S3,EN_REGR=>EN_REGR_S3,ENABLE=>ENABLE_S3,SEL2=> SEL2_S3,EN_REGO=>EN_REGO_S3,WR=>P_7,WI=>N_7, CLK=>CLK,SEL_INV=>SEL_INV_S3);
BF_3_3: BF PORT MAP(AI=>S23_2_BI,AR=>S23_2_BR,BR=>S23_3_BR,BI=>S23_3_BI, A1R=>C3AR_OUT,A1I=>C3AI_OUT,B1R=>							C3BR_OUT,B1I=>C3BI_OUT,SEL3=>SEL3_S3,SEL1=>SEL1_S3,SELSUM=>SELSUM_S3,C=>C_S3,A_S=>							A_S_S3,EN_REGR=>EN_REGR_S3,ENABLE=>ENABLE_S3,SEL2=> SEL2_S3,EN_REGO=>EN_REGO_S3,WR=>N_7,WI=>N_7, CLK=>CLK,SEL_INV=>SEL_INV_S3);
BF_3_4: BF PORT MAP(AI=>S23_4_AI,AR=>S23_4_AR,BR=>S23_5_AR,BI=>S23_5_AI, A1R=>C4AR_OUT,A1I=>C4AI_OUT,B1R=>							C4BR_OUT,B1I=>C4BI_OUT,SEL3=>SEL3_S3,SEL1=>SEL1_S3,SELSUM=>SELSUM_S3,C=>C_S3,A_S=>							A_S_S3,EN_REGR=>EN_REGR_S3,ENABLE=>ENABLE_S3,SEL2=> SEL2_S3,EN_REGO=>EN_REGO_S3,WR=>P_9,WI=>N_3, CLK=>CLK,SEL_INV=>SEL_INV_S3);
BF_3_5: BF PORT MAP(AI=>S23_4_BI,AR=>S23_4_BR,BR=>S23_5_BR,BI=>S23_5_BI, A1R=>C5AR_OUT,A1I=>C5AI_OUT,B1R=>							C5BR_OUT,B1I=>C5BI_OUT,SEL3=>SEL3_S3,SEL1=>SEL1_S3,SELSUM=>SELSUM_S3,C=>C_S3,A_S=>							A_S_S3,EN_REGR=>EN_REGR_S3,ENABLE=>ENABLE_S3,SEL2=> SEL2_S3,EN_REGO=>EN_REGO_S3,WR=>N_3,WI=>N_9, CLK=>CLK,SEL_INV=>SEL_INV_S3);
BF_3_6: BF PORT MAP(AI=>S23_6_AI,AR=>S23_6_AR,BR=>S23_7_AR,BI=>S23_7_AI, A1R=>C6AR_OUT,A1I=>C6AI_OUT,B1R=>							C6BR_OUT,B1I=>C6BI_OUT,SEL3=>SEL3_S3,SEL1=>SEL1_S3,SELSUM=>SELSUM_S3,C=>C_S3,A_S=>							A_S_S3,EN_REGR=>EN_REGR_S3,ENABLE=>ENABLE_S3,SEL2=> SEL2_S3,EN_REGO=>EN_REGO_S3,WR=>P_3,WI=>N_9, CLK=>CLK,SEL_INV=>SEL_INV_S3);
BF_3_7: BF PORT MAP(AI=>S23_6_BI,AR=>S23_6_BR,BR=>S23_7_BR,BI=>S23_7_BI, A1R=>C7AR_OUT,A1I=>C7AI_OUT,B1R=>							C7BR_OUT,B1I=>C7BI_OUT,SEL3=>SEL3_S3,SEL1=>SEL1_S3,SELSUM=>SELSUM_S3,C=>C_S3,A_S=>							A_S_S3,EN_REGR=>EN_REGR_S3,ENABLE=>ENABLE_S3,SEL2=> SEL2_S3,EN_REGO=>EN_REGO_S3,WR=>N_9,WI=>N_3, CLK=>CLK,SEL_INV=>SEL_INV_S3);

OR_LOGIC:OR_PORT PORT MAP(START=>START_S,B0AR=>C0AR,B1AR=>C1AR,B2AR=>C2AR,B3AR=>C3AR,B4AR=>C4AR,B5AR=>C5AR,									B6AR=>C6AR,B7AR=>C7AR,
								 B0AI=>C0AI,B1AI=>C1AI,B2AI=>C2AI,B3AI=>C3AI,B4AI=>C4AI,B5AI=>C5AI,B6AI=>C6AI,B7AI								  =>C7AI,B0BR=>C0BR,B1BR=>C1BR,B2BR=>C2BR,B3BR=>C3BR,B4BR=>C4BR,B5BR=>C5BR,B6BR=>								 C6BR,B7BR=>C7BR,B0BI=>C0BI,B1BI=>C1BI,B2BI=>C2BI,B3BI=>C3BI,B4BI=>C4BI,B5BI=>C5BI,								   B6BI=>C6BI,B7BI=>C7BI);
								 
								 
SEQ_LOGIC: XOR_CHECK PORT MAP(OUT_XOR_CHECK=>OUT_XOR_CHECK_S,B0AR=>C0AR_GUARD_S,B1AR=>C1AR_GUARD_S,B2AR=>C2AR_GUARD_S,B3AR=>C3AR_GUARD_S,								B4AR=>C4AR_GUARD_S,B5AR=>C5AR_GUARD_S,B6AR=>C6AR_GUARD_S,B7AR=>C7AR_GUARD_S,B0AI=>C0AI_GUARD_S,B1AI=>C1AI_GUARD_S,B2AI=>C2AI_GUARD_S,B3AI=>								C3AI_GUARD_S,B4AI=>C4AI_GUARD_S,B5AI=>C5AI_GUARD_S,B6AI=>C6AI_GUARD_S,B7AI=>C7AI_GUARD_S,B0BR=>C0BR_GUARD_S,B1BR=>C1BR_GUARD_S,B2BR=>C2BR_GUARD_S,							 B3BR=>C3BR_GUARD_S,B4BR=>C4BR_GUARD_S,B5BR=>C5BR_GUARD_S,B6BR=>C6BR_GUARD_S,B7BR=>C7BR_GUARD_S,B0BI=>C0BI_GUARD_S,B1BI=>C1BI_GUARD_S,B2BI=>							C2BI_GUARD_S,B3BI=>C3BI_GUARD_S,B4BI=>C4BI_GUARD_S,B5BI=>C5BI_GUARD_S,B6BI=>C6BI_GUARD_S,B7BI=>C7BI_GUARD_S,B0AR_OLD=>AR0_CTRL,								B1AR_OLD=>AR1_CTRL,B2AR_OLD=>AR2_CTRL,B3AR_OLD=>AR3_CTRL,B4AR_OLD=>AR4_CTRL,							B5AR_OLD=>AR5_CTRL,B6AR_OLD=>AR6_CTRL,B7AR_OLD=>AR7_CTRL,B0AI_OLD=>AI0_CTRL,B1AI_OLD=>							AI1_CTRL,B2AI_OLD=>AI2_CTRL,B3AI_OLD=>AI3_CTRL,B4AI_OLD=>AI4_CTRL,B5AI_OLD=>AI5_CTRL,							B6AI_OLD=>AI6_CTRL,B7AI_OLD=>AI7_CTRL,B0BR_OLD=>BR0_CTRL,B1BR_OLD=>BR1_CTRL,B2BR_OLD=>							BR2_CTRL,B3BR_OLD=>BR3_CTRL,B4BR_OLD=>BR4_CTRL,B5BR_OLD=>BR5_CTRL,B6BR_OLD=>BR6_CTRL,							B7BR_OLD=>BR7_CTRL,B0BI_OLD=>BI0_CTRL,B1BI_OLD=>BI1_CTRL,B2BI_OLD=>BI2_CTRL,B3BI_OLD=>							BI3_CTRL,B4BI_OLD=>BI4_CTRL,B5BI_OLD=>BI5_CTRL,B6BI_OLD=>BI6_CTRL,B7BI_OLD=>BI7_CTRL);	

STONE_0:	R_STONE_0 PORT MAP(OUTPUT=>P_0);				 
STONE_1: R_STONE_1 PORT MAP(OUTPUT_P=>P_1,OUTPUT_N=>N_1);	
STONE_3: R_STONE_3 PORT MAP(OUTPUT_P=>P_3,OUTPUT_N=>N_3);
STONE_7: R_STONE_7 PORT MAP(OUTPUT_P=>P_7,OUTPUT_N=>N_7);
STONE_9: R_STONE_9 PORT MAP(OUTPUT_P=>P_9,OUTPUT_N=>N_9);

-- CU BF
CU0 : CU_BF PORT MAP (LOAD=>ENABLE_S0,SEQ=>SEQ_CU0,CLK=>CLK,RESET=>RESET,CTRL_OUT(14)=>SEL_INV_S0,
							 CTRL_OUT(13)=>SELSUM_S0,CTRL_OUT(12)=>SEL1_S0,CTRL_OUT(11 downto 10)=>SEL2_S0,
							 CTRL_OUT(9)=>SEL3_S0,CTRL_OUT(8)=>C_S0,CTRL_OUT(7)=>A_S_S0,CTRL_OUT(6)=>EN_REGS0,
							 CTRL_OUT(5)=>EN_REGR_S0,CTRL_OUT(4 DOWNTO 2)=>EN_REGO_S0,CTRL_OUT(1)=>FREE_M_TOP,
							 CTRL_OUT(0)=>ENABLE_S1);
CU1 : CU_BF PORT MAP (LOAD=>ENABLE_S1,SEQ=>SEQ_CU1,CLK=>CLK,RESET=>RESET,CTRL_OUT(14)=>SEL_INV_S1,
							 CTRL_OUT(13)=>SELSUM_S1,CTRL_OUT(12)=>SEL1_S1,CTRL_OUT(11 downto 10)=>SEL2_S1,
							 CTRL_OUT(9)=>SEL3_S1,CTRL_OUT(8)=>C_S1,CTRL_OUT(7)=>A_S_S1,CTRL_OUT(6)=>EN_REGS1,
							 CTRL_OUT(5)=>EN_REGR_S1,CTRL_OUT(4 DOWNTO 2)=>EN_REGO_S1,CTRL_OUT(1)=>FREE_M_S,
							 CTRL_OUT(0)=>ENABLE_S2);
CU2 : CU_BF PORT MAP (LOAD=>ENABLE_S2,SEQ=>SEQ_CU2,CLK=>CLK,RESET=>RESET,CTRL_OUT(14)=>SEL_INV_S2,
							 CTRL_OUT(13)=>SELSUM_S2,CTRL_OUT(12)=>SEL1_S2,CTRL_OUT(11 downto 10)=>SEL2_S2,
							 CTRL_OUT(9)=>SEL3_S2,CTRL_OUT(8)=>C_S2,CTRL_OUT(7)=>A_S_S2,CTRL_OUT(6)=>EN_REGS2,
							 CTRL_OUT(5)=>EN_REGR_S2,CTRL_OUT(4 DOWNTO 2)=>EN_REGO_S2,CTRL_OUT(1)=>FREE_M_S,
							 CTRL_OUT(0)=>ENABLE_S3);
CU3 : CU_BF PORT MAP (LOAD=>ENABLE_S3,SEQ=>SEQ_CU3,CLK=>CLK,RESET=>RESET,CTRL_OUT(14)=>SEL_INV_S3,
							 CTRL_OUT(13)=>SELSUM_S3,CTRL_OUT(12)=>SEL1_S3,CTRL_OUT(11 downto 10)=>SEL2_S3,
							 CTRL_OUT(9)=>SEL3_S3,CTRL_OUT(8)=>C_S3,CTRL_OUT(7)=>A_S_S3,CTRL_OUT(6)=>EN_REGS3,
							 CTRL_OUT(5)=>EN_REGR_S3,CTRL_OUT(4 DOWNTO 2)=>EN_REGO_S3,CTRL_OUT(1)=>FREE_M_S,
							 CTRL_OUT(0)=>END_BF_TOP);

--CU TOP
TOP : CU_TOP PORT MAP (START=>START_S_TOP,PROGRESS=>NEW_PROGRESS_S,FREE_M=>FREE_M_TOP,END_BF=>END_BF_TOP,
							  SEQ=>NEW_OUT_XOR_CHECK_S,CLK=>CLK,RESET=>RESET,
							  CTRL_TOP_OUT(5)=>ENABLE_S0,CTRL_TOP_OUT(4)=>EN_FF_S,CTRL_TOP_OUT(3)=>FF_VALUE_S,
							  CTRL_TOP_OUT(2)=>DONE,CTRL_TOP_OUT(1)=>READY,CTRL_TOP_OUT(0)=>RESET_OUT);
							  
-- SENSE START
SS : start_sense PORT MAP(D=>EN_FF_S,CLK=>CLK,set=>RESET_OUT,enable=>EN_FF_S,SENSE=>SENSE_S);

-- REG STATUS
RS : REG_STATUS PORT MAP (CLK=>CLK,set=>ENABLE_S0,enable0=>EN_REGS0,enable1=>EN_REGS1,enable2=>EN_REGS2,
								  enable3=>EN_REGS3,Q_OUT=>PROGRESS_S,RESET=>RESET_OUT);
-- REG SEQ
RSEQ : REG_SEQ PORT MAP (CLK=>CLK,D0=>NEW_OUT_XOR_CHECK_S,D1=>PROGRESS_S(0),D2=>PROGRESS_S(1),D3=>PROGRESS_S(2),
								 SET=>SET_REG_SEQ,RESET=>RESET_OUT,EN0=>ENABLE_S1,EN1=>ENABLE_S2,
						EN2=>ENABLE_S3,EN3=>END_BF_TOP,Q0=>SEQ_CU0,Q1=>SEQ_CU1,Q2=>SEQ_CU2,Q3=>SEQ_CU3);

GB : GUARD PORT MAP (C0AR=>C0AR,C1AR=>C1AR,C2AR=>C2AR,C3AR=>C3AR,C4AR=>C4AR,C5AR=>C5AR,C6AR=>C6AR,C7AR=>C7AR,
							C0AI=>C0AI,C1AI=>C1AI,C2AI=>C2AI,C3AI=>C3AI,C4AI=>C4AI,C5AI=>C5AI,C6AI=>C6AI,C7AI=>C7AI,
							C0BR=>C0BR,C1BR=>C1BR,C2BR=>C2BR,C3BR=>C3BR,C4BR=>C4BR,C5BR=>C5BR,C6BR=>C6BR,C7BR=>C7BR,
							C0BI=>C0BI,C1BI=>C1BI,C2BI=>C2BI,C3BI=>C3BI,C4BI=>C4BI,C5BI=>C5BI,C6BI=>C6BI,C7BI=>C7BI,
							
							C0AR_GUARD=>C0AR_GUARD_S,C1AR_GUARD=>C1AR_GUARD_S,C2AR_GUARD=>C2AR_GUARD_S,C3AR_GUARD=>C3AR_GUARD_S,
							C4AR_GUARD=>C4AR_GUARD_S,C5AR_GUARD=>C5AR_GUARD_S,C6AR_GUARD=>C6AR_GUARD_S,C7AR_GUARD=>C7AR_GUARD_S,
							C0AI_GUARD=>C0AI_GUARD_S,C1AI_GUARD=>C1AI_GUARD_S,C2AI_GUARD=>C2AI_GUARD_S,C3AI_GUARD=>C3AI_GUARD_S,
							C4AI_GUARD=>C4AI_GUARD_S,C5AI_GUARD=>C5AI_GUARD_S,C6AI_GUARD=>C6AI_GUARD_S,C7AI_GUARD=>C7AI_GUARD_S, 
							C0BR_GUARD=>C0BR_GUARD_S,C1BR_GUARD=>C1BR_GUARD_S,C2BR_GUARD=>C2BR_GUARD_S,C3BR_GUARD=>C3BR_GUARD_S,
							C4BR_GUARD=>C4BR_GUARD_S,C5BR_GUARD=>C5BR_GUARD_S,C6BR_GUARD=>C6BR_GUARD_S,C7BR_GUARD=>C7BR_GUARD_S, 
							C0BI_GUARD=>C0BI_GUARD_S,C1BI_GUARD=>C1BI_GUARD_S,C2BI_GUARD=>C2BI_GUARD_S,C3BI_GUARD=>C3BI_GUARD_S,
							C4BI_GUARD=>C4BI_GUARD_S,C5BI_GUARD=>C5BI_GUARD_S,C6BI_GUARD=>C6BI_GUARD_S,C7BI_GUARD=>C7BI_GUARD_S); 							 	
	
END BEHAV;