LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all; 

ENTITY R_STONE_7 IS

PORT(
      OUTPUT_P,OUTPUT_N: OUT SIGNED(19 DOWNTO 0));
END R_STONE_7;


ARCHITECTURE BEHAV OF R_STONE_7 IS 
SIGNAL VALORE :SIGNED (19 DOWNTO 0);
BEGIN  --
--VALORE<= "01011010100000000000";
VALORE<= "01011010100000101000";
OUTPUT_P<=VALORE;
OUTPUT_N(19 downto 4)<= NOT VALORE(19 downto 4);
OUTPUT_N(3 downto 0)<= VALORE(3 DOWNTO 0);
END BEHAV;