LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all; 


ENTITY FFT_16_tb IS 
END FFT_16_tb;

ARCHITECTURE behav OF FFT_16_tb IS

SIGNAL CLK_tb,RESET_tb,DONE_tb,READY_tb:STD_LOGIC;
SIGNAL C0AR_tb,C1AR_tb,C2AR_tb,C3AR_tb,C4AR_tb,C5AR_tb,C6AR_tb,C7AR_tb: SIGNED(19 downto 0);
SIGNAL C0AI_tb,C1AI_tb,C2AI_tb,C3AI_tb,C4AI_tb,C5AI_tb,C6AI_tb,C7AI_tb: SIGNED(19 downto 0);
SIGNAL C0BR_tb,C1BR_tb,C2BR_tb,C3BR_tb,C4BR_tb,C5BR_tb,C6BR_tb,C7BR_tb: SIGNED(19 downto 0);
SIGNAL C0BI_tb,C1BI_tb,C2BI_tb,C3BI_tb,C4BI_tb,C5BI_tb,C6BI_tb,C7BI_tb: SIGNED(19 downto 0);
		
SIGNAL C0AR_OUT_tb,C1AR_OUT_tb,C2AR_OUT_tb,C3AR_OUT_tb,C4AR_OUT_tb,C5AR_OUT_tb,C6AR_OUT_tb,C7AR_OUT_tb: SIGNED(19 downto 0);
SIGNAL C0AI_OUT_tb,C1AI_OUT_tb,C2AI_OUT_tb,C3AI_OUT_tb,C4AI_OUT_tb,C5AI_OUT_tb,C6AI_OUT_tb,C7AI_OUT_tb: SIGNED(19 downto 0);
SIGNAL C0BR_OUT_tb,C1BR_OUT_tb,C2BR_OUT_tb,C3BR_OUT_tb,C4BR_OUT_tb,C5BR_OUT_tb,C6BR_OUT_tb,C7BR_OUT_tb: SIGNED(19 downto 0);
SIGNAL C0BI_OUT_tb,C1BI_OUT_tb,C2BI_OUT_tb,C3BI_OUT_tb,C4BI_OUT_tb,C5BI_OUT_tb,C6BI_OUT_tb,C7BI_OUT_tb: SIGNED(19 downto 0);


COMPONENT FFT_16 IS
PORT ( CLK,RESET: IN STD_LOGIC;
		 DONE,READY: OUT STD_LOGIC;
       C0AR,C1AR,C2AR,C3AR,C4AR,C5AR,C6AR,C7AR: IN SIGNED(19 downto 0);
		 C0AI,C1AI,C2AI,C3AI,C4AI,C5AI,C6AI,C7AI: IN SIGNED(19 downto 0);
		 C0BR,C1BR,C2BR,C3BR,C4BR,C5BR,C6BR,C7BR: IN SIGNED(19 downto 0);
		 C0BI,C1BI,C2BI,C3BI,C4BI,C5BI,C6BI,C7BI: IN SIGNED(19 downto 0);
		
	    C0AR_OUT,C1AR_OUT,C2AR_OUT,C3AR_OUT,C4AR_OUT,C5AR_OUT,C6AR_OUT,C7AR_OUT: 
		 OUT SIGNED(19 downto 0);
		 C0AI_OUT,C1AI_OUT,C2AI_OUT,C3AI_OUT,C4AI_OUT,C5AI_OUT,C6AI_OUT,C7AI_OUT: 
		 OUT SIGNED(19 downto 0);
		 C0BR_OUT,C1BR_OUT,C2BR_OUT,C3BR_OUT,C4BR_OUT,C5BR_OUT,C6BR_OUT,C7BR_OUT: 
		 OUT SIGNED(19 downto 0);
		 C0BI_OUT,C1BI_OUT,C2BI_OUT,C3BI_OUT,C4BI_OUT,C5BI_OUT,C6BI_OUT,C7BI_OUT: 
		 OUT SIGNED(19 downto 0));
END COMPONENT;

BEGIN

FFT: FFT_16 PORT MAP(CLK=>CLK_tb,RESET=>RESET_tb,DONE=>DONE_tb,READY=>READY_tb,

C0AR=>C0AR_tb,C1AR=>C1AR_tb,C2AR=>C2AR_tb,C3AR=>C3AR_tb,C4AR=>C4AR_tb,C5AR=>C5AR_tb,C6AR=>C6AR_tb,C7AR=>C7AR_tb,
C0AI=>C0AI_tb,C1AI=>C1AI_tb,C2AI=>C2AI_tb,C3AI=>C3AI_tb,C4AI=>C4AI_tb,C5AI=>C5AI_tb,C6AI=>C6AI_tb,C7AI=>C7AI_tb,
C0BR=>C0BR_tb,C1BR=>C1BR_tb,C2BR=>C2BR_tb,C3BR=>C3BR_tb,C4BR=>C4BR_tb,C5BR=>C5BR_tb,C6BR=>C6BR_tb,C7BR=>C7BR_tb,
C0BI=>C0BI_tb,C1BI=>C1BI_tb,C2BI=>C2BI_tb,C3BI=>C3BI_tb,C4BI=>C4BI_tb,C5BI=>C5BI_tb,C6BI=>C6BI_tb,C7BI=>C7BI_tb,

							C0AR_OUT=>C0AR_OUT_tb,C1AR_OUT=>C1AR_OUT_tb,C2AR_OUT=>C2AR_OUT_tb,C3AR_OUT=>C3AR_OUT_tb,
							C4AR_OUT=>C4AR_OUT_tb,C5AR_OUT=>C5AR_OUT_tb,C6AR_OUT=>C6AR_OUT_tb,C7AR_OUT=>C7AR_OUT_tb,
							
							C0AI_OUT=>C0AI_OUT_tb,C1AI_OUT=>C1AI_OUT_tb,C2AI_OUT=>C2AI_OUT_tb,C3AI_OUT=>C3AI_OUT_tb,
							C4AI_OUT=>C4AI_OUT_tb,C5AI_OUT=>C5AI_OUT_tb,C6AI_OUT=>C6AI_OUT_tb,C7AI_OUT=>C7AI_OUT_tb,
							
							C0BR_OUT=>C0BR_OUT_tb,C1BR_OUT=>C1BR_OUT_tb,C2BR_OUT=>C2BR_OUT_tb,C3BR_OUT=>C3BR_OUT_tb,
							C4BR_OUT=>C4BR_OUT_tb,C5BR_OUT=>C5BR_OUT_tb,C6BR_OUT=>C6BR_OUT_tb,C7BR_OUT=>C7BR_OUT_tb,
							
							C0BI_OUT=>C0BI_OUT_tb,C1BI_OUT=>C1BI_OUT_tb,C2BI_OUT=>C2BI_OUT_tb,C3BI_OUT=>C3BI_OUT_tb,
							C4BI_OUT=>C4BI_OUT_tb,C5BI_OUT=>C5BI_OUT_tb,C6BI_OUT=>C6BI_OUT_tb,C7BI_OUT=>C7BI_OUT_tb);
							
 clk_process: PROCESS 
 
 BEGIN 
 CLK_tb<= '0';
 wait for 10 ns;	
 CLK_tb <= '1';
 wait for 10 ns;
 end process;
 
 --  0 : 00000000000000000000
 -- -1 : 10000000000000000000
 --  1 : 01111111111111111111
 -- 0.5: 01000000000000000000
 -- -0.5:11000000000000000000
 -- 0.75:01100000000000000000
 
 ingressi: PROCESS
 BEGIN
 C0AR_tb<="00000000000000000000"; 
 C1AR_tb<="00000000000000000000"; 
 C2AR_tb<="00000000000000000000";
 C3AR_tb<="00000000000000000000";
 C4AR_tb<="00000000000000000000";
 C5AR_tb<="00000000000000000000";
 C6AR_tb<="00000000000000000000";
 C7AR_tb<="00000000000000000000";
 C0AI_tb<="00000000000000000000";
 C1AI_tb<="00000000000000000000";
 C2AI_tb<="00000000000000000000";
 C3AI_tb<="00000000000000000000";
 C4AI_tb<="00000000000000000000";
 C5AI_tb<="00000000000000000000";
 C6AI_tb<="00000000000000000000";
 C7AI_tb<="00000000000000000000";
 C0BR_tb<="00000000000000000000";
 C1BR_tb<="00000000000000000000";
 C2BR_tb<="00000000000000000000";
 C3BR_tb<="00000000000000000000";
 C4BR_tb<="00000000000000000000";
 C5BR_tb<="00000000000000000000";
 C6BR_tb<="00000000000000000000";
 C7BR_tb<="00000000000000000000";
 C0BI_tb<="00000000000000000000";
 C1BI_tb<="00000000000000000000";
 C2BI_tb<="00000000000000000000";
 C3BI_tb<="00000000000000000000";
 C4BI_tb<="00000000000000000000";
 C5BI_tb<="00000000000000000000";
 C6BI_tb<="00000000000000000000";
 C7BI_tb<="00000000000000000000";
 wait for 50 ns;
 -- CAMPIONE 1
 C0AR_tb<="10000000000000000000"; 
 C1AR_tb<="10000000000000000000"; 
 C2AR_tb<="10000000000000000000";
 C3AR_tb<="10000000000000000000";
 C4AR_tb<="10000000000000000000";
 C5AR_tb<="10000000000000000000";
 C6AR_tb<="10000000000000000000";
 C7AR_tb<="10000000000000000000";
 C0AI_tb<="00000000000000000000";
 C1AI_tb<="00000000000000000000";
 C2AI_tb<="00000000000000000000";
 C3AI_tb<="00000000000000000000";
 C4AI_tb<="00000000000000000000";
 C5AI_tb<="00000000000000000000";
 C6AI_tb<="00000000000000000000";
 C7AI_tb<="00000000000000000000";
 C0BR_tb<="10000000000000000000";
 C1BR_tb<="10000000000000000000";
 C2BR_tb<="10000000000000000000";
 C3BR_tb<="10000000000000000000";
 C4BR_tb<="10000000000000000000";
 C5BR_tb<="10000000000000000000";
 C6BR_tb<="10000000000000000000";
 C7BR_tb<="10000000000000000000";
 C0BI_tb<="00000000000000000000";
 C1BI_tb<="00000000000000000000";
 C2BI_tb<="00000000000000000000";
 C3BI_tb<="00000000000000000000";
 C4BI_tb<="00000000000000000000";
 C5BI_tb<="00000000000000000000";
 C6BI_tb<="00000000000000000000";
 C7BI_tb<="00000000000000000000";
 wait for 140 ns;
 -- CAMPIONE 2
 C0AR_tb<="10000000000000000000"; 
C1AR_tb<="00000000000000000000"; 
C2AR_tb<="01111111111111111111";
C3AR_tb<="00000000000000000000";
C4AR_tb<="10000000000000000000";
C5AR_tb<="00000000000000000000";
C6AR_tb<="01111111111111111111";
C7AR_tb<="00000000000000000000";
C0AI_tb<="00000000000000000000";
C1AI_tb<="00000000000000000000";
C2AI_tb<="00000000000000000000";
C3AI_tb<="00000000000000000000";
C4AI_tb<="00000000000000000000";
C5AI_tb<="00000000000000000000";
C6AI_tb<="00000000000000000000";
C7AI_tb<="00000000000000000000";
C0BR_tb<="10000000000000000000";
C1BR_tb<="00000000000000000000";
C2BR_tb<="01111111111111111111";
C3BR_tb<="00000000000000000000";
C4BR_tb<="10000000000000000000";
C5BR_tb<="00000000000000000000";
C6BR_tb<="01111111111111111111";
C7BR_tb<="00000000000000000000";
C0BI_tb<="00000000000000000000";
C1BI_tb<="00000000000000000000";
C2BI_tb<="00000000000000000000";
C3BI_tb<="00000000000000000000";
C4BI_tb<="00000000000000000000";
C5BI_tb<="00000000000000000000";
C6BI_tb<="00000000000000000000";
C7BI_tb<="00000000000000000000";
 wait for 140 ns;
 -- CAMPIONE 3
 C0AR_tb<="01111111111111111111"; 
 C1AR_tb<="00000000000000000000"; 
 C2AR_tb<="00000000000000000000";
 C3AR_tb<="00000000000000000000";
 C4AR_tb<="00000000000000000000";
 C5AR_tb<="00000000000000000000";
 C6AR_tb<="00000000000000000000";
 C7AR_tb<="00000000000000000000";
 C0AI_tb<="00000000000000000000";
 C1AI_tb<="00000000000000000000";
 C2AI_tb<="00000000000000000000";
 C3AI_tb<="00000000000000000000";
 C4AI_tb<="00000000000000000000";
 C5AI_tb<="00000000000000000000";
 C6AI_tb<="00000000000000000000";
 C7AI_tb<="00000000000000000000";
 C0BR_tb<="00000000000000000000";
 C1BR_tb<="00000000000000000000";
 C2BR_tb<="00000000000000000000";
 C3BR_tb<="00000000000000000000";
 C4BR_tb<="00000000000000000000";
 C5BR_tb<="00000000000000000000";
 C6BR_tb<="00000000000000000000";
 C7BR_tb<="00000000000000000000";
 C0BI_tb<="00000000000000000000";
 C1BI_tb<="00000000000000000000";
 C2BI_tb<="00000000000000000000";
 C3BI_tb<="00000000000000000000";
 C4BI_tb<="00000000000000000000";
 C5BI_tb<="00000000000000000000";
 C6BI_tb<="00000000000000000000";
 C7BI_tb<="00000000000000000000";
 wait for 140 ns;
 -- CAMPIONE 4
 C0AR_tb<="10000000000000000000"; 
 C1AR_tb<="10000000000000000000"; 
 C2AR_tb<="01111111111111111111";
 C3AR_tb<="01111111111111111111";
 C4AR_tb<="10000000000000000000";
 C5AR_tb<="10000000000000000000";
 C6AR_tb<="01111111111111111111";
 C7AR_tb<="01111111111111111111";
 C0AI_tb<="00000000000000000000";
 C1AI_tb<="00000000000000000000";
 C2AI_tb<="00000000000000000000";
 C3AI_tb<="00000000000000000000";
 C4AI_tb<="00000000000000000000";
 C5AI_tb<="00000000000000000000";
 C6AI_tb<="00000000000000000000";
 C7AI_tb<="00000000000000000000";
 C0BR_tb<="10000000000000000000";
 C1BR_tb<="10000000000000000000";
 C2BR_tb<="01111111111111111111";
 C3BR_tb<="01111111111111111111";
 C4BR_tb<="10000000000000000000";
 C5BR_tb<="10000000000000000000";
 C6BR_tb<="01111111111111111111";
 C7BR_tb<="01111111111111111111";
 C0BI_tb<="00000000000000000000";
 C1BI_tb<="00000000000000000000";
 C2BI_tb<="00000000000000000000";
 C3BI_tb<="00000000000000000000";
 C4BI_tb<="00000000000000000000";
 C5BI_tb<="00000000000000000000";
 C6BI_tb<="00000000000000000000";
 C7BI_tb<="00000000000000000000";
 wait for 140 ns;
 -- CAMPIONE 5
 C0AR_tb<="01000000000000000000"; 
 C1AR_tb<="01000000000000000000"; 
 C2AR_tb<="01000000000000000000";
 C3AR_tb<="01000000000000000000";
 C4AR_tb<="01000000000000000000";
 C5AR_tb<="01000000000000000000";
 C6AR_tb<="01000000000000000000";
 C7AR_tb<="01000000000000000000";
 C0AI_tb<="00000000000000000000";
 C1AI_tb<="00000000000000000000";
 C2AI_tb<="00000000000000000000";
 C3AI_tb<="00000000000000000000";
 C4AI_tb<="00000000000000000000";
 C5AI_tb<="00000000000000000000";
 C6AI_tb<="00000000000000000000";
 C7AI_tb<="00000000000000000000";
 C0BR_tb<="01000000000000000000";
 C1BR_tb<="11000000000000000000";
 C2BR_tb<="11000000000000000000";
 C3BR_tb<="11000000000000000000";
 C4BR_tb<="11000000000000000000";
 C5BR_tb<="11000000000000000000";
 C6BR_tb<="11000000000000000000";
 C7BR_tb<="11000000000000000000";
 C0BI_tb<="00000000000000000000";
 C1BI_tb<="00000000000000000000";
 C2BI_tb<="00000000000000000000";
 C3BI_tb<="00000000000000000000";
 C4BI_tb<="00000000000000000000";
 C5BI_tb<="00000000000000000000";
 C6BI_tb<="00000000000000000000";
 C7BI_tb<="00000000000000000000";
 wait for 140 ns;
 -- CAMPIONE 6
 C0AR_tb<="00000000000000000000"; 
 C1AR_tb<="00000000000000000000"; 
 C2AR_tb<="00000000000000000000";
 C3AR_tb<="00000000000000000000";
 C4AR_tb<="00000000000000000000";
 C5AR_tb<="00000000000000000000";
 C6AR_tb<="00000000000000000000";
 C7AR_tb<="00000000000000000000";
 C0AI_tb<="00000000000000000000";
 C1AI_tb<="00000000000000000000";
 C2AI_tb<="00000000000000000000";
 C3AI_tb<="00000000000000000000";
 C4AI_tb<="00000000000000000000";
 C5AI_tb<="00000000000000000000";
 C6AI_tb<="00000000000000000000";
 C7AI_tb<="00000000000000000000";
 C0BR_tb<="01100000000000000000";
 C1BR_tb<="00000000000000000000";
 C2BR_tb<="00000000000000000000";
 C3BR_tb<="00000000000000000000";
 C4BR_tb<="00000000000000000000";
 C5BR_tb<="00000000000000000000";
 C6BR_tb<="00000000000000000000";
 C7BR_tb<="00000000000000000000";
 C0BI_tb<="00000000000000000000";
 C1BI_tb<="00000000000000000000";
 C2BI_tb<="00000000000000000000";
 C3BI_tb<="00000000000000000000";
 C4BI_tb<="00000000000000000000";
 C5BI_tb<="00000000000000000000";
 C6BI_tb<="00000000000000000000";
 C7BI_tb<="00000000000000000000";
 wait for 140 ns;
 C0AR_tb<="00000000000000000000"; 
 C1AR_tb<="00000000000000000000"; 
 C2AR_tb<="00000000000000000000";
 C3AR_tb<="00000000000000000000";
 C4AR_tb<="00000000000000000000";
 C5AR_tb<="00000000000000000000";
 C6AR_tb<="00000000000000000000";
 C7AR_tb<="00000000000000000000";
 C0AI_tb<="00000000000000000000";
 C1AI_tb<="00000000000000000000";
 C2AI_tb<="00000000000000000000";
 C3AI_tb<="00000000000000000000";
 C4AI_tb<="00000000000000000000";
 C5AI_tb<="00000000000000000000";
 C6AI_tb<="00000000000000000000";
 C7AI_tb<="00000000000000000000";
 C0BR_tb<="00000000000000000000";
 C1BR_tb<="00000000000000000000";
 C2BR_tb<="00000000000000000000";
 C3BR_tb<="00000000000000000000";
 C4BR_tb<="00000000000000000000";
 C5BR_tb<="00000000000000000000";
 C6BR_tb<="00000000000000000000";
 C7BR_tb<="00000000000000000000";
 C0BI_tb<="00000000000000000000";
 C1BI_tb<="00000000000000000000";
 C2BI_tb<="00000000000000000000";
 C3BI_tb<="00000000000000000000";
 C4BI_tb<="00000000000000000000";
 C5BI_tb<="00000000000000000000";
 C6BI_tb<="00000000000000000000";
 C7BI_tb<="00000000000000000000";
 wait for 5000 ns;
 END PROCESS;
 
 PROCESS
 BEGIN
 RESET_tb<='1';
 wait for 10 ns;
 RESET_tb<='0';
 wait for 10000 ns;
 END PROCESS;
 END behav;