LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all; 

ENTITY R_STONE_3 IS

PORT(
      OUTPUT_P,OUTPUT_N: OUT SIGNED(19 DOWNTO 0));
END R_STONE_3;


ARCHITECTURE BEHAV OF R_STONE_3 IS 
SIGNAL VALORE :SIGNED (19 DOWNTO 0);
BEGIN  
--VALORE<= "00110000111100000000";
VALORE<= "00110000111110111100";
OUTPUT_P<=VALORE;
OUTPUT_N(19 downto 3)<= NOT VALORE(19 downto 3);
OUTPUT_N(2 downto 0)<= VALORE(2 DOWNTO 0);
END BEHAV;